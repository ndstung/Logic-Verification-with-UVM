// output is real, imag
// real is rv[45:23]
// imag is rv[22:0]
function reg [45:0] fftwiddle(reg [5:0] ix);
    reg [45:0] rv;
    case(ix)
      0 : rv={23'd32768, 23'd0};
      1 : rv={23'd32728, -23'd1607};
      2 : rv={23'd32610, -23'd3211};
      3 : rv={23'd32413, -23'd4808};
      4 : rv={23'd32138, -23'd6392};
      5 : rv={23'd31785, -23'd7961};
      6 : rv={23'd31357, -23'd9512};
      7 : rv={23'd30852, -23'd11039};
      8 : rv={23'd30273, -23'd12539};
      9 : rv={23'd29621, -23'd14010};
      10 : rv={23'd28898, -23'd15446};
      11 : rv={23'd28106, -23'd16846};
      12 : rv={23'd27245, -23'd18204};
      13 : rv={23'd26319, -23'd19519};
      14 : rv={23'd25330, -23'd20787};
      15 : rv={23'd24279, -23'd22005};
      16 : rv={23'd23170, -23'd23170};
      17 : rv={23'd22005, -23'd24279};
      18 : rv={23'd20787, -23'd25330};
      19 : rv={23'd19519, -23'd26319};
      20 : rv={23'd18204, -23'd27245};
      21 : rv={23'd16846, -23'd28106};
      22 : rv={23'd15446, -23'd28898};
      23 : rv={23'd14010, -23'd29621};
      24 : rv={23'd12539, -23'd30273};
      25 : rv={23'd11039, -23'd30852};
      26 : rv={23'd9512, -23'd31357};
      27 : rv={23'd7961, -23'd31785};
      28 : rv={23'd6392, -23'd32138};
      29 : rv={23'd4808, -23'd32413};
      30 : rv={23'd3211, -23'd32610};
      31 : rv={23'd1607, -23'd32728};
      32 : rv={23'd0, -23'd32768};
      33 : rv={-23'd1607, -23'd32728};
      34 : rv={-23'd3211, -23'd32610};
      35 : rv={-23'd4808, -23'd32413};
      36 : rv={-23'd6392, -23'd32138};
      37 : rv={-23'd7961, -23'd31785};
      38 : rv={-23'd9512, -23'd31357};
      39 : rv={-23'd11039, -23'd30852};
      40 : rv={-23'd12539, -23'd30273};
      41 : rv={-23'd14010, -23'd29621};
      42 : rv={-23'd15446, -23'd28898};
      43 : rv={-23'd16846, -23'd28106};
      44 : rv={-23'd18204, -23'd27245};
      45 : rv={-23'd19519, -23'd26319};
      46 : rv={-23'd20787, -23'd25330};
      47 : rv={-23'd22005, -23'd24279};
      48 : rv={-23'd23170, -23'd23170};
      49 : rv={-23'd24279, -23'd22005};
      50 : rv={-23'd25330, -23'd20787};
      51 : rv={-23'd26319, -23'd19519};
      52 : rv={-23'd27245, -23'd18204};
      53 : rv={-23'd28106, -23'd16846};
      54 : rv={-23'd28898, -23'd15446};
      55 : rv={-23'd29621, -23'd14010};
      56 : rv={-23'd30273, -23'd12539};
      57 : rv={-23'd30852, -23'd11039};
      58 : rv={-23'd31357, -23'd9512};
      59 : rv={-23'd31785, -23'd7961};
      60 : rv={-23'd32138, -23'd6392};
      61 : rv={-23'd32413, -23'd4808};
      62 : rv={-23'd32610, -23'd3211};
      63 : rv={-23'd32728, -23'd1607};
    endcase
    return rv;
  endfunction : fftwiddle
  